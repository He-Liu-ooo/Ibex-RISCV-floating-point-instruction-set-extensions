module sram_32x1024
(
  input  logic       CLK,
  input  logic       RSTN,
  input  logic       CEN,
  input  logic       WEN,
  input  logic [9:0] A,
  input  logic [31:0] D,
  output logic [31:0] Q
);

  logic [31:0] mem [1023:0];

  always_ff @(posedge CLK or negedge RSTN) begin
    if(!RSTN) begin
      // 17
      mem[0] = 32'h0;
      mem[1] = 32'h3F400000;
      mem[2] = 32'h42960000;
      mem[3] = 32'h42700000;
      mem[4] = 32'h42E60000;
      mem[5] = 32'h42BE0000;
      mem[6] = 32'h0;
      mem[7] = 32'h1;
      mem[8] = 32'h1;
      mem[9] = 32'h3F68F5C2;
      mem[10] = 32'h42A00000;
      mem[11] = 32'h42700000;
      mem[12] = 32'h42F00000;
      mem[13] = 32'h42C80000;
      mem[14] = 32'h0;
      mem[15] = 32'h1;
      mem[16] = 32'h2;
      mem[17] = 32'h3F23D70A;
      mem[18] = 32'h42AA0000;
      mem[19] = 32'h42820000;
      mem[20] = 32'h42FA0000;
      mem[21] = 32'h42D20000;
      mem[22] = 32'h0;
      mem[23] = 32'h1;
      mem[24] = 32'h3;
      mem[25] = 32'h3F333333;
      mem[26] = 32'h42B40000;
      mem[27] = 32'h425C0000;
      mem[28] = 32'h42FA0000;
      mem[29] = 32'h42C80000;
      mem[30] = 32'h0;
      mem[31] = 32'h1;
      mem[32] = 32'h4;
      mem[33] = 32'h3F63D70A;
      mem[34] = 32'h41700000;
      mem[35] = 32'h42BE0000;
      mem[36] = 32'h420C0000;
      mem[37] = 32'h42F00000;
      mem[38] = 32'h0;
      mem[39] = 32'h1;
      mem[40] = 32'h5;
      mem[41] = 32'h3F4A3D70;
      mem[42] = 32'h41200000;
      mem[43] = 32'h42B40000;
      mem[44] = 32'h41F00000;
      mem[45] = 32'h42E60000;
      mem[46] = 32'h0;
      mem[47] = 32'h1;
      mem[48] = 32'h6;
      mem[49] = 32'h3F35C28F;
      mem[50] = 32'h431B0000;
      mem[51] = 32'h42C80000;
      mem[52] = 32'h43390000;
      mem[53] = 32'h43020000;
      mem[54] = 32'h0;
      mem[55] = 32'h1;
      mem[56] = 32'h7;
      mem[57] = 32'h3F63D70A;
      mem[58] = 32'h43250000;
      mem[59] = 32'h42BE0000;
      mem[60] = 32'h433E0000;
      mem[61] = 32'h43070000;
      mem[62] = 32'h0;
      mem[63] = 32'h1;
      mem[64] = 32'h8;
      mem[65] = 32'h3F68F5C2;
      mem[66] = 32'h43200000;
      mem[67] = 32'h42D20000;
      mem[68] = 32'h433E0000;
      mem[69] = 32'h42FA0000;
      mem[70] = 32'h0;
      mem[71] = 32'h1;
      mem[72] = 32'h9;
      mem[73] = 32'h3F547AE1;
      mem[74] = 32'h41A00000;
      mem[75] = 32'h41A00000;
      mem[76] = 32'h42820000;
      mem[77] = 32'h42960000;
      mem[78] = 32'h1;
      mem[79] = 32'h1;
      mem[80] = 32'ha;
      mem[81] = 32'h3F400000;
      mem[82] = 32'h40A00000;
      mem[83] = 32'h41700000;
      mem[84] = 32'h425C0000;
      mem[85] = 32'h42820000;
      mem[86] = 32'h1;
      mem[87] = 32'h1;
      mem[88] = 32'hb;
      mem[89] = 32'h3F7AE147;
      mem[90] = 32'h41200000;
      mem[91] = 32'h41A00000;
      mem[92] = 32'h42700000;
      mem[93] = 32'h428C0000;
      mem[94] = 32'h1;
      mem[95] = 32'h1;
      mem[96] = 32'hc;
      mem[97] = 32'h3F2B851E;
      mem[98] = 32'h431B0000;
      mem[99] = 32'h420C0000;
      mem[100] = 32'h434D0000;
      mem[101] = 32'h42AA0000;
      mem[102] = 32'h2;
      mem[103] = 32'h1;
      mem[104] = 32'hd;
      mem[105] = 32'h3F4F5C28;
      mem[106] = 32'h43160000;
      mem[107] = 32'h41F00000;
      mem[108] = 32'h43480000;
      mem[109] = 32'h42A00000;
      mem[110] = 32'h2;
      mem[111] = 32'h1;
      mem[112] = 32'he;
      mem[113] = 32'h3F5EB851;
      mem[114] = 32'h42B40000;
      mem[115] = 32'h41200000;
      mem[116] = 32'h42F00000;
      mem[117] = 32'h42200000;
      mem[118] = 32'h2;
      mem[119] = 32'h1;
      mem[120] = 32'hf;
      mem[121] = 32'h3F666666;
      mem[122] = 32'h42C80000;
      mem[123] = 32'h41200000;
      mem[124] = 32'h42FA0000;
      mem[125] = 32'h420C0000;
      mem[126] = 32'h2;
      mem[127] = 32'h1;
      mem[128] = 32'h10;
      mem[129] = 32'h3F599999;
      mem[130] = 32'h42BE0000;
      mem[131] = 32'h40A00000;
      mem[132] = 32'h42F00000;
      mem[133] = 32'h41F00000;
      mem[134] = 32'h2;
      mem[135] = 32'h1;

      // 14
      //       mem[0] = 32'h0;
//       mem[1] = 32'h3fe00000;
//       mem[2] = 32'h40a00000;
//       mem[3] = 32'h40a00000;
//       mem[4] = 32'h425c0000;
//       mem[5] = 32'h428c0000;
//       mem[6] = 32'h0;
//       mem[7] = 32'h1;
//       mem[8] = 32'h1;
//       mem[9] = 32'h3fea3d70;
//       mem[10] = 32'h41200000;
//       mem[11] = 32'h41200000;
//       mem[12] = 32'h42700000;
//       mem[13] = 32'h42960000;
//       mem[14] = 32'h0;
//       mem[15] = 32'h1;
//       mem[16] = 32'h2;
//       mem[17] = 32'h3fdae147;
//       mem[18] = 32'h41700000;
//       mem[19] = 32'h40a00000;
//       mem[20] = 32'h428c0000;
//       mem[21] = 32'h42820000;
//       mem[22] = 32'h0;
//       mem[23] = 32'h1;
//       mem[24] = 32'h3;
//       mem[25] = 32'h3FE7AE14;
//       mem[26] = 32'h42820000;
//       mem[27] = 32'h42BE0000;
//       mem[28] = 32'h42C80000;
//       mem[29] = 32'h430C0000;
//       mem[30] = 32'h0;
//       mem[31] = 32'h1;
//       mem[32] = 32'h4;
//       mem[33] = 32'h3FFC28F5;
//       mem[34] = 32'h428C0000;
//       mem[35] = 32'h42C80000;
//       mem[36] = 32'h42BE0000;
//       mem[37] = 32'h43070000;
//       mem[38] = 32'h0;
//       mem[39] = 32'h1;
//       mem[40] = 32'h5;
//       mem[41] = 32'h3FE51EB8;
//       mem[42] = 32'h42B40000;
//       mem[43] = 32'h42820000;
//       mem[44] = 32'h42FA0000;
//       mem[45] = 32'h42D20000;
//       mem[46] = 32'h1;
//       mem[47] = 32'h1;
//       mem[48] = 32'h6;
//       mem[49] = 32'h3FE7AE14;
//       mem[50] = 32'h42BE0000;
//       mem[51] = 32'h428C0000;
//       mem[52] = 32'h43020000;
//       mem[53] = 32'h42DC0000;
//       mem[54] = 32'h1;
//       mem[55] = 32'h1;
//       mem[56] = 32'h7;
//       mem[57] = 32'h3FF5C28F;
//       mem[58] = 32'h42C80000;
//       mem[59] = 32'h42820000;
//       mem[60] = 32'h43020000;
//       mem[61] = 32'h42E60000;
//       mem[62] = 32'h1;
//       mem[63] = 32'h1;
//       mem[64] = 32'h8;
//       mem[65] = 32'h3ff33333;
//       mem[66] = 32'h41200000;
//       mem[67] = 32'h42be0000;
//       mem[68] = 32'h420c0000;
//       mem[69] = 32'h42f00000;
//       mem[70] = 32'h1;
//       mem[71] = 32'h1;
//       mem[72] = 32'h9;
//       mem[73] = 32'h3fe66666;
//       mem[74] = 32'h41700000;
//       mem[75] = 32'h42aa0000;
//       mem[76] = 32'h42200000;
//       mem[77] = 32'h42e60000;
//       mem[78] = 32'h1;
//       mem[79] = 32'h1;
//       mem[80] = 32'ha;
//       mem[81] = 32'h3FEF5C28;
//       mem[82] = 32'h43020000;
//       mem[83] = 32'h40A00000;
//       mem[84] = 32'h43340000;
//       mem[85] = 32'h42340000;
//       mem[86] = 32'h1;
//       mem[87] = 32'h1;
//       mem[88] = 32'hb;
//       mem[89] = 32'h3FF47AE1;
//       mem[90] = 32'h43070000;
//       mem[91] = 32'h00000000;
//       mem[92] = 32'h43390000;
//       mem[93] = 32'h42480000;
//       mem[94] = 32'h1;
//       mem[95] = 32'h1;
//       mem[96] = 32'hc;
//       mem[97] = 32'h3FF99999;
//       mem[98] = 32'h430C0000;
//       mem[99] = 32'h40A00000;
//       mem[100] = 32'h43340000;
//       mem[101] = 32'h425C0000;
//       mem[102] = 32'h1;
//       mem[103] = 32'h1;
//       mem[104] = 32'hd;
//       mem[105] = 32'h3FE147AE;
//       mem[106] = 32'h43110000;
//       mem[107] = 32'h41200000;
//       mem[108] = 32'h43390000;
//       mem[109] = 32'h42700000;
//       mem[110] = 32'h1;
//       mem[111] = 32'h1;
      
    end 
    else if(!CEN&&!WEN)  // 两者同为低的时候才能写入
      mem[A] <= D;
    else ;
  end

  always_ff@(posedge CLK) begin
    if(!CEN&&WEN)     // CEN 为低，写使能为高的时候才能读出
      Q <= mem[A];
  end
  
endmodule

